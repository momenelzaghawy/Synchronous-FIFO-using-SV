package internal_pkg;
bit test_finished ;
integer error_count=0,correct_count=0;
    
endpackage